module erl

fn C.enif_get_int(&u8, DynamicTerm, &u8) int