module erl

fn C.enif_make_string(&u8, &u8, Encoding) DynamicTerm
fn C.enif_make_int(&u8, int) DynamicTerm
fn C.enif_make_badarg(&u8) DynamicTerm